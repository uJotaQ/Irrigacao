module main();
	
endmodule
