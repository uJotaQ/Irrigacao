module Aspersao(AS, GT_wire, US);
	input GT_wire, US;
	output AS;
	
	nor NotOr0(AS, GT_wire, US);
	
endmodule